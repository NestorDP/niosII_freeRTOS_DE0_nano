// niosII.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module niosII (
		input  wire        clk_clk,            //         clk.clk
		output wire        epcs_dclk,          //        epcs.dclk
		output wire        epcs_sce,           //            .sce
		output wire        epcs_sdo,           //            .sdo
		input  wire        epcs_data0,         //            .data0
		inout  wire [31:0] port_gpio_0_export, // port_gpio_0.export
		input  wire [1:0]  port_key_export,    //    port_key.export
		output wire [7:0]  port_led_export,    //    port_led.export
		input  wire [3:0]  port_sw_export,     //     port_sw.export
		output wire        ram_clk_clk,        //     ram_clk.clk
		input  wire        reset_reset_n,      //       reset.reset_n
		output wire [12:0] sdram_addr,         //       sdram.addr
		output wire [1:0]  sdram_ba,           //            .ba
		output wire        sdram_cas_n,        //            .cas_n
		output wire        sdram_cke,          //            .cke
		output wire        sdram_cs_n,         //            .cs_n
		inout  wire [15:0] sdram_dq,           //            .dq
		output wire [1:0]  sdram_dqm,          //            .dqm
		output wire        sdram_ras_n,        //            .ras_n
		output wire        sdram_we_n,         //            .we_n
		input  wire        uart_rxd,           //        uart.rxd
		output wire        uart_txd            //            .txd
	);

	wire         sys_pll_c0_clk;                                                     // sys_pll:c0 -> [Button_Pio:clk, IO_Pio:clk, LED_Pio:clk, Switch_Pio:clk, cpu:clk, epcs:clk, irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:receiver_clk, irq_synchronizer_001:sender_clk, mm_interconnect_0:sys_clk_clk_clk, mm_interconnect_0:sys_pll_c0_clk, rst_controller:clk, rst_controller_001:clk, sdram:clk, sys_clk_timer:clk, sys_id:clock, uart:clk]
	wire  [31:0] cpu_data_master_readdata;                                           // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                                        // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                                        // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [26:0] cpu_data_master_address;                                            // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                         // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                               // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_write;                                              // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                          // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                                    // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                                 // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [26:0] cpu_instruction_master_address;                                     // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                        // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;                // mm_interconnect_0:jtag_avalon_jtag_slave_chipselect -> jtag:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;                  // jtag:av_readdata -> mm_interconnect_0:jtag_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest;               // jtag:av_waitrequest -> mm_interconnect_0:jtag_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;                   // mm_interconnect_0:jtag_avalon_jtag_slave_address -> jtag:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;                      // mm_interconnect_0:jtag_avalon_jtag_slave_read -> jtag:av_read_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;                     // mm_interconnect_0:jtag_avalon_jtag_slave_write -> jtag:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;                 // mm_interconnect_0:jtag_avalon_jtag_slave_writedata -> jtag:av_writedata
	wire         mm_interconnect_0_led_pio_avalon_parallel_port_slave_chipselect;    // mm_interconnect_0:LED_Pio_avalon_parallel_port_slave_chipselect -> LED_Pio:chipselect
	wire  [31:0] mm_interconnect_0_led_pio_avalon_parallel_port_slave_readdata;      // LED_Pio:readdata -> mm_interconnect_0:LED_Pio_avalon_parallel_port_slave_readdata
	wire   [1:0] mm_interconnect_0_led_pio_avalon_parallel_port_slave_address;       // mm_interconnect_0:LED_Pio_avalon_parallel_port_slave_address -> LED_Pio:address
	wire         mm_interconnect_0_led_pio_avalon_parallel_port_slave_read;          // mm_interconnect_0:LED_Pio_avalon_parallel_port_slave_read -> LED_Pio:read
	wire   [3:0] mm_interconnect_0_led_pio_avalon_parallel_port_slave_byteenable;    // mm_interconnect_0:LED_Pio_avalon_parallel_port_slave_byteenable -> LED_Pio:byteenable
	wire         mm_interconnect_0_led_pio_avalon_parallel_port_slave_write;         // mm_interconnect_0:LED_Pio_avalon_parallel_port_slave_write -> LED_Pio:write
	wire  [31:0] mm_interconnect_0_led_pio_avalon_parallel_port_slave_writedata;     // mm_interconnect_0:LED_Pio_avalon_parallel_port_slave_writedata -> LED_Pio:writedata
	wire         mm_interconnect_0_button_pio_avalon_parallel_port_slave_chipselect; // mm_interconnect_0:Button_Pio_avalon_parallel_port_slave_chipselect -> Button_Pio:chipselect
	wire  [31:0] mm_interconnect_0_button_pio_avalon_parallel_port_slave_readdata;   // Button_Pio:readdata -> mm_interconnect_0:Button_Pio_avalon_parallel_port_slave_readdata
	wire   [1:0] mm_interconnect_0_button_pio_avalon_parallel_port_slave_address;    // mm_interconnect_0:Button_Pio_avalon_parallel_port_slave_address -> Button_Pio:address
	wire         mm_interconnect_0_button_pio_avalon_parallel_port_slave_read;       // mm_interconnect_0:Button_Pio_avalon_parallel_port_slave_read -> Button_Pio:read
	wire   [3:0] mm_interconnect_0_button_pio_avalon_parallel_port_slave_byteenable; // mm_interconnect_0:Button_Pio_avalon_parallel_port_slave_byteenable -> Button_Pio:byteenable
	wire         mm_interconnect_0_button_pio_avalon_parallel_port_slave_write;      // mm_interconnect_0:Button_Pio_avalon_parallel_port_slave_write -> Button_Pio:write
	wire  [31:0] mm_interconnect_0_button_pio_avalon_parallel_port_slave_writedata;  // mm_interconnect_0:Button_Pio_avalon_parallel_port_slave_writedata -> Button_Pio:writedata
	wire         mm_interconnect_0_switch_pio_avalon_parallel_port_slave_chipselect; // mm_interconnect_0:Switch_Pio_avalon_parallel_port_slave_chipselect -> Switch_Pio:chipselect
	wire  [31:0] mm_interconnect_0_switch_pio_avalon_parallel_port_slave_readdata;   // Switch_Pio:readdata -> mm_interconnect_0:Switch_Pio_avalon_parallel_port_slave_readdata
	wire   [1:0] mm_interconnect_0_switch_pio_avalon_parallel_port_slave_address;    // mm_interconnect_0:Switch_Pio_avalon_parallel_port_slave_address -> Switch_Pio:address
	wire         mm_interconnect_0_switch_pio_avalon_parallel_port_slave_read;       // mm_interconnect_0:Switch_Pio_avalon_parallel_port_slave_read -> Switch_Pio:read
	wire   [3:0] mm_interconnect_0_switch_pio_avalon_parallel_port_slave_byteenable; // mm_interconnect_0:Switch_Pio_avalon_parallel_port_slave_byteenable -> Switch_Pio:byteenable
	wire         mm_interconnect_0_switch_pio_avalon_parallel_port_slave_write;      // mm_interconnect_0:Switch_Pio_avalon_parallel_port_slave_write -> Switch_Pio:write
	wire  [31:0] mm_interconnect_0_switch_pio_avalon_parallel_port_slave_writedata;  // mm_interconnect_0:Switch_Pio_avalon_parallel_port_slave_writedata -> Switch_Pio:writedata
	wire         mm_interconnect_0_io_pio_avalon_parallel_port_slave_chipselect;     // mm_interconnect_0:IO_Pio_avalon_parallel_port_slave_chipselect -> IO_Pio:chipselect
	wire  [31:0] mm_interconnect_0_io_pio_avalon_parallel_port_slave_readdata;       // IO_Pio:readdata -> mm_interconnect_0:IO_Pio_avalon_parallel_port_slave_readdata
	wire   [1:0] mm_interconnect_0_io_pio_avalon_parallel_port_slave_address;        // mm_interconnect_0:IO_Pio_avalon_parallel_port_slave_address -> IO_Pio:address
	wire         mm_interconnect_0_io_pio_avalon_parallel_port_slave_read;           // mm_interconnect_0:IO_Pio_avalon_parallel_port_slave_read -> IO_Pio:read
	wire   [3:0] mm_interconnect_0_io_pio_avalon_parallel_port_slave_byteenable;     // mm_interconnect_0:IO_Pio_avalon_parallel_port_slave_byteenable -> IO_Pio:byteenable
	wire         mm_interconnect_0_io_pio_avalon_parallel_port_slave_write;          // mm_interconnect_0:IO_Pio_avalon_parallel_port_slave_write -> IO_Pio:write
	wire  [31:0] mm_interconnect_0_io_pio_avalon_parallel_port_slave_writedata;      // mm_interconnect_0:IO_Pio_avalon_parallel_port_slave_writedata -> IO_Pio:writedata
	wire  [31:0] mm_interconnect_0_sys_id_control_slave_readdata;                    // sys_id:readdata -> mm_interconnect_0:sys_id_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sys_id_control_slave_address;                     // mm_interconnect_0:sys_id_control_slave_address -> sys_id:address
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;                     // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;                  // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;                  // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;                      // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                         // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;                   // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;                        // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;                    // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire         mm_interconnect_0_epcs_epcs_control_port_chipselect;                // mm_interconnect_0:epcs_epcs_control_port_chipselect -> epcs:chipselect
	wire  [31:0] mm_interconnect_0_epcs_epcs_control_port_readdata;                  // epcs:readdata -> mm_interconnect_0:epcs_epcs_control_port_readdata
	wire   [8:0] mm_interconnect_0_epcs_epcs_control_port_address;                   // mm_interconnect_0:epcs_epcs_control_port_address -> epcs:address
	wire         mm_interconnect_0_epcs_epcs_control_port_read;                      // mm_interconnect_0:epcs_epcs_control_port_read -> epcs:read_n
	wire         mm_interconnect_0_epcs_epcs_control_port_write;                     // mm_interconnect_0:epcs_epcs_control_port_write -> epcs:write_n
	wire  [31:0] mm_interconnect_0_epcs_epcs_control_port_writedata;                 // mm_interconnect_0:epcs_epcs_control_port_writedata -> epcs:writedata
	wire  [31:0] mm_interconnect_0_sys_pll_pll_slave_readdata;                       // sys_pll:readdata -> mm_interconnect_0:sys_pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_sys_pll_pll_slave_address;                        // mm_interconnect_0:sys_pll_pll_slave_address -> sys_pll:address
	wire         mm_interconnect_0_sys_pll_pll_slave_read;                           // mm_interconnect_0:sys_pll_pll_slave_read -> sys_pll:read
	wire         mm_interconnect_0_sys_pll_pll_slave_write;                          // mm_interconnect_0:sys_pll_pll_slave_write -> sys_pll:write
	wire  [31:0] mm_interconnect_0_sys_pll_pll_slave_writedata;                      // mm_interconnect_0:sys_pll_pll_slave_writedata -> sys_pll:writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                              // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                                // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                             // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [23:0] mm_interconnect_0_sdram_s1_address;                                 // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                    // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                              // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                           // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                   // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                               // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_sys_clk_timer_s1_chipselect;                      // mm_interconnect_0:sys_clk_timer_s1_chipselect -> sys_clk_timer:chipselect
	wire  [15:0] mm_interconnect_0_sys_clk_timer_s1_readdata;                        // sys_clk_timer:readdata -> mm_interconnect_0:sys_clk_timer_s1_readdata
	wire   [2:0] mm_interconnect_0_sys_clk_timer_s1_address;                         // mm_interconnect_0:sys_clk_timer_s1_address -> sys_clk_timer:address
	wire         mm_interconnect_0_sys_clk_timer_s1_write;                           // mm_interconnect_0:sys_clk_timer_s1_write -> sys_clk_timer:write_n
	wire  [15:0] mm_interconnect_0_sys_clk_timer_s1_writedata;                       // mm_interconnect_0:sys_clk_timer_s1_writedata -> sys_clk_timer:writedata
	wire         mm_interconnect_0_uart_s1_chipselect;                               // mm_interconnect_0:uart_s1_chipselect -> uart:chipselect
	wire  [15:0] mm_interconnect_0_uart_s1_readdata;                                 // uart:readdata -> mm_interconnect_0:uart_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_s1_address;                                  // mm_interconnect_0:uart_s1_address -> uart:address
	wire         mm_interconnect_0_uart_s1_read;                                     // mm_interconnect_0:uart_s1_read -> uart:read_n
	wire         mm_interconnect_0_uart_s1_begintransfer;                            // mm_interconnect_0:uart_s1_begintransfer -> uart:begintransfer
	wire         mm_interconnect_0_uart_s1_write;                                    // mm_interconnect_0:uart_s1_write -> uart:write_n
	wire  [15:0] mm_interconnect_0_uart_s1_writedata;                                // mm_interconnect_0:uart_s1_writedata -> uart:writedata
	wire         irq_mapper_receiver1_irq;                                           // sys_clk_timer:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver3_irq;                                           // uart:irq -> irq_mapper:receiver3_irq
	wire  [31:0] cpu_irq_irq;                                                        // irq_mapper:sender_irq -> cpu:irq
	wire         irq_mapper_receiver0_irq;                                           // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                      // jtag:av_irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver2_irq;                                           // irq_synchronizer_001:sender_irq -> irq_mapper:receiver2_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                                  // epcs:irq -> irq_synchronizer_001:receiver_irq
	wire         rst_controller_reset_out_reset;                                     // rst_controller:reset_out -> [Button_Pio:reset, IO_Pio:reset, LED_Pio:reset, Switch_Pio:reset, cpu:reset_n, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, sdram:reset_n, sys_clk_timer:reset_n, sys_id:reset_n, uart:reset_n]
	wire         rst_controller_reset_out_reset_req;                                 // rst_controller:reset_req -> [cpu:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                                 // rst_controller_001:reset_out -> [epcs:reset_n, irq_synchronizer_001:receiver_reset, mm_interconnect_0:epcs_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset_req;                             // rst_controller_001:reset_req -> [epcs:reset_req, rst_translator_001:reset_req_in]
	wire         cpu_debug_reset_request_reset;                                      // cpu:debug_reset_request -> rst_controller_001:reset_in1
	wire         rst_controller_002_reset_out_reset;                                 // rst_controller_002:reset_out -> [irq_synchronizer:receiver_reset, jtag:rst_n, mm_interconnect_0:jtag_reset_reset_bridge_in_reset_reset, sys_pll:reset]

	niosII_Button_Pio button_pio (
		.clk        (sys_pll_c0_clk),                                                     //                        clk.clk
		.reset      (rst_controller_reset_out_reset),                                     //                      reset.reset
		.address    (mm_interconnect_0_button_pio_avalon_parallel_port_slave_address),    // avalon_parallel_port_slave.address
		.byteenable (mm_interconnect_0_button_pio_avalon_parallel_port_slave_byteenable), //                           .byteenable
		.chipselect (mm_interconnect_0_button_pio_avalon_parallel_port_slave_chipselect), //                           .chipselect
		.read       (mm_interconnect_0_button_pio_avalon_parallel_port_slave_read),       //                           .read
		.write      (mm_interconnect_0_button_pio_avalon_parallel_port_slave_write),      //                           .write
		.writedata  (mm_interconnect_0_button_pio_avalon_parallel_port_slave_writedata),  //                           .writedata
		.readdata   (mm_interconnect_0_button_pio_avalon_parallel_port_slave_readdata),   //                           .readdata
		.KEY        (port_key_export)                                                     //         external_interface.export
	);

	niosII_IO_Pio io_pio (
		.clk        (sys_pll_c0_clk),                                                 //                        clk.clk
		.reset      (rst_controller_reset_out_reset),                                 //                      reset.reset
		.address    (mm_interconnect_0_io_pio_avalon_parallel_port_slave_address),    // avalon_parallel_port_slave.address
		.byteenable (mm_interconnect_0_io_pio_avalon_parallel_port_slave_byteenable), //                           .byteenable
		.chipselect (mm_interconnect_0_io_pio_avalon_parallel_port_slave_chipselect), //                           .chipselect
		.read       (mm_interconnect_0_io_pio_avalon_parallel_port_slave_read),       //                           .read
		.write      (mm_interconnect_0_io_pio_avalon_parallel_port_slave_write),      //                           .write
		.writedata  (mm_interconnect_0_io_pio_avalon_parallel_port_slave_writedata),  //                           .writedata
		.readdata   (mm_interconnect_0_io_pio_avalon_parallel_port_slave_readdata),   //                           .readdata
		.GPIO_0     (port_gpio_0_export)                                              //         external_interface.export
	);

	niosII_LED_Pio led_pio (
		.clk        (sys_pll_c0_clk),                                                  //                        clk.clk
		.reset      (rst_controller_reset_out_reset),                                  //                      reset.reset
		.address    (mm_interconnect_0_led_pio_avalon_parallel_port_slave_address),    // avalon_parallel_port_slave.address
		.byteenable (mm_interconnect_0_led_pio_avalon_parallel_port_slave_byteenable), //                           .byteenable
		.chipselect (mm_interconnect_0_led_pio_avalon_parallel_port_slave_chipselect), //                           .chipselect
		.read       (mm_interconnect_0_led_pio_avalon_parallel_port_slave_read),       //                           .read
		.write      (mm_interconnect_0_led_pio_avalon_parallel_port_slave_write),      //                           .write
		.writedata  (mm_interconnect_0_led_pio_avalon_parallel_port_slave_writedata),  //                           .writedata
		.readdata   (mm_interconnect_0_led_pio_avalon_parallel_port_slave_readdata),   //                           .readdata
		.LEDG       (port_led_export)                                                  //         external_interface.export
	);

	niosII_Switch_Pio switch_pio (
		.clk        (sys_pll_c0_clk),                                                     //                        clk.clk
		.reset      (rst_controller_reset_out_reset),                                     //                      reset.reset
		.address    (mm_interconnect_0_switch_pio_avalon_parallel_port_slave_address),    // avalon_parallel_port_slave.address
		.byteenable (mm_interconnect_0_switch_pio_avalon_parallel_port_slave_byteenable), //                           .byteenable
		.chipselect (mm_interconnect_0_switch_pio_avalon_parallel_port_slave_chipselect), //                           .chipselect
		.read       (mm_interconnect_0_switch_pio_avalon_parallel_port_slave_read),       //                           .read
		.write      (mm_interconnect_0_switch_pio_avalon_parallel_port_slave_write),      //                           .write
		.writedata  (mm_interconnect_0_switch_pio_avalon_parallel_port_slave_writedata),  //                           .writedata
		.readdata   (mm_interconnect_0_switch_pio_avalon_parallel_port_slave_readdata),   //                           .readdata
		.DIP        (port_sw_export)                                                      //         external_interface.export
	);

	niosII_cpu cpu (
		.clk                                 (sys_pll_c0_clk),                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	niosII_epcs epcs (
		.clk        (sys_pll_c0_clk),                                      //               clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                 //             reset.reset_n
		.reset_req  (rst_controller_001_reset_out_reset_req),              //                  .reset_req
		.address    (mm_interconnect_0_epcs_epcs_control_port_address),    // epcs_control_port.address
		.chipselect (mm_interconnect_0_epcs_epcs_control_port_chipselect), //                  .chipselect
		.read_n     (~mm_interconnect_0_epcs_epcs_control_port_read),      //                  .read_n
		.readdata   (mm_interconnect_0_epcs_epcs_control_port_readdata),   //                  .readdata
		.write_n    (~mm_interconnect_0_epcs_epcs_control_port_write),     //                  .write_n
		.writedata  (mm_interconnect_0_epcs_epcs_control_port_writedata),  //                  .writedata
		.irq        (irq_synchronizer_001_receiver_irq),                   //               irq.irq
		.dclk       (epcs_dclk),                                           //          external.export
		.sce        (epcs_sce),                                            //                  .export
		.sdo        (epcs_sdo),                                            //                  .export
		.data0      (epcs_data0)                                           //                  .export
	);

	niosII_jtag jtag (
		.clk            (clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                  //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_synchronizer_receiver_irq)                         //               irq.irq
	);

	niosII_sdram sdram (
		.clk            (sys_pll_c0_clk),                           //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	niosII_sys_clk_timer sys_clk_timer (
		.clk        (sys_pll_c0_clk),                                //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               // reset.reset_n
		.address    (mm_interconnect_0_sys_clk_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_sys_clk_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_sys_clk_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_sys_clk_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_sys_clk_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                       //   irq.irq
	);

	niosII_sys_id sys_id (
		.clock    (sys_pll_c0_clk),                                  //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                 //         reset.reset_n
		.readdata (mm_interconnect_0_sys_id_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sys_id_control_slave_address)   //              .address
	);

	niosII_sys_pll sys_pll (
		.clk                (clk_clk),                                       //       inclk_interface.clk
		.reset              (rst_controller_002_reset_out_reset),            // inclk_interface_reset.reset
		.read               (mm_interconnect_0_sys_pll_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_sys_pll_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_sys_pll_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_sys_pll_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_sys_pll_pll_slave_writedata), //                      .writedata
		.c0                 (sys_pll_c0_clk),                                //                    c0.clk
		.c1                 (ram_clk_clk),                                   //                    c1.clk
		.scandone           (),                                              //           (terminated)
		.scandataout        (),                                              //           (terminated)
		.areset             (1'b0),                                          //           (terminated)
		.locked             (),                                              //           (terminated)
		.phasedone          (),                                              //           (terminated)
		.phasecounterselect (4'b0000),                                       //           (terminated)
		.phaseupdown        (1'b0),                                          //           (terminated)
		.phasestep          (1'b0),                                          //           (terminated)
		.scanclk            (1'b0),                                          //           (terminated)
		.scanclkena         (1'b0),                                          //           (terminated)
		.scandata           (1'b0),                                          //           (terminated)
		.configupdate       (1'b0)                                           //           (terminated)
	);

	niosII_uart uart (
		.clk           (sys_pll_c0_clk),                          //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address       (mm_interconnect_0_uart_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_s1_readdata),      //                    .readdata
		.rxd           (uart_rxd),                                // external_connection.export
		.txd           (uart_txd),                                //                    .export
		.irq           (irq_mapper_receiver3_irq)                 //                 irq.irq
	);

	niosII_mm_interconnect_0 mm_interconnect_0 (
		.clock_50_clk_clk                                 (clk_clk),                                                            //                          clock_50_clk.clk
		.sys_clk_clk_clk                                  (sys_pll_c0_clk),                                                     //                           sys_clk_clk.clk
		.sys_pll_c0_clk                                   (sys_pll_c0_clk),                                                     //                            sys_pll_c0.clk
		.cpu_reset_reset_bridge_in_reset_reset            (rst_controller_reset_out_reset),                                     //       cpu_reset_reset_bridge_in_reset.reset
		.epcs_reset_reset_bridge_in_reset_reset           (rst_controller_001_reset_out_reset),                                 //      epcs_reset_reset_bridge_in_reset.reset
		.jtag_reset_reset_bridge_in_reset_reset           (rst_controller_002_reset_out_reset),                                 //      jtag_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                          (cpu_data_master_address),                                            //                       cpu_data_master.address
		.cpu_data_master_waitrequest                      (cpu_data_master_waitrequest),                                        //                                      .waitrequest
		.cpu_data_master_byteenable                       (cpu_data_master_byteenable),                                         //                                      .byteenable
		.cpu_data_master_read                             (cpu_data_master_read),                                               //                                      .read
		.cpu_data_master_readdata                         (cpu_data_master_readdata),                                           //                                      .readdata
		.cpu_data_master_write                            (cpu_data_master_write),                                              //                                      .write
		.cpu_data_master_writedata                        (cpu_data_master_writedata),                                          //                                      .writedata
		.cpu_data_master_debugaccess                      (cpu_data_master_debugaccess),                                        //                                      .debugaccess
		.cpu_instruction_master_address                   (cpu_instruction_master_address),                                     //                cpu_instruction_master.address
		.cpu_instruction_master_waitrequest               (cpu_instruction_master_waitrequest),                                 //                                      .waitrequest
		.cpu_instruction_master_read                      (cpu_instruction_master_read),                                        //                                      .read
		.cpu_instruction_master_readdata                  (cpu_instruction_master_readdata),                                    //                                      .readdata
		.Button_Pio_avalon_parallel_port_slave_address    (mm_interconnect_0_button_pio_avalon_parallel_port_slave_address),    // Button_Pio_avalon_parallel_port_slave.address
		.Button_Pio_avalon_parallel_port_slave_write      (mm_interconnect_0_button_pio_avalon_parallel_port_slave_write),      //                                      .write
		.Button_Pio_avalon_parallel_port_slave_read       (mm_interconnect_0_button_pio_avalon_parallel_port_slave_read),       //                                      .read
		.Button_Pio_avalon_parallel_port_slave_readdata   (mm_interconnect_0_button_pio_avalon_parallel_port_slave_readdata),   //                                      .readdata
		.Button_Pio_avalon_parallel_port_slave_writedata  (mm_interconnect_0_button_pio_avalon_parallel_port_slave_writedata),  //                                      .writedata
		.Button_Pio_avalon_parallel_port_slave_byteenable (mm_interconnect_0_button_pio_avalon_parallel_port_slave_byteenable), //                                      .byteenable
		.Button_Pio_avalon_parallel_port_slave_chipselect (mm_interconnect_0_button_pio_avalon_parallel_port_slave_chipselect), //                                      .chipselect
		.cpu_debug_mem_slave_address                      (mm_interconnect_0_cpu_debug_mem_slave_address),                      //                   cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                        (mm_interconnect_0_cpu_debug_mem_slave_write),                        //                                      .write
		.cpu_debug_mem_slave_read                         (mm_interconnect_0_cpu_debug_mem_slave_read),                         //                                      .read
		.cpu_debug_mem_slave_readdata                     (mm_interconnect_0_cpu_debug_mem_slave_readdata),                     //                                      .readdata
		.cpu_debug_mem_slave_writedata                    (mm_interconnect_0_cpu_debug_mem_slave_writedata),                    //                                      .writedata
		.cpu_debug_mem_slave_byteenable                   (mm_interconnect_0_cpu_debug_mem_slave_byteenable),                   //                                      .byteenable
		.cpu_debug_mem_slave_waitrequest                  (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),                  //                                      .waitrequest
		.cpu_debug_mem_slave_debugaccess                  (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),                  //                                      .debugaccess
		.epcs_epcs_control_port_address                   (mm_interconnect_0_epcs_epcs_control_port_address),                   //                epcs_epcs_control_port.address
		.epcs_epcs_control_port_write                     (mm_interconnect_0_epcs_epcs_control_port_write),                     //                                      .write
		.epcs_epcs_control_port_read                      (mm_interconnect_0_epcs_epcs_control_port_read),                      //                                      .read
		.epcs_epcs_control_port_readdata                  (mm_interconnect_0_epcs_epcs_control_port_readdata),                  //                                      .readdata
		.epcs_epcs_control_port_writedata                 (mm_interconnect_0_epcs_epcs_control_port_writedata),                 //                                      .writedata
		.epcs_epcs_control_port_chipselect                (mm_interconnect_0_epcs_epcs_control_port_chipselect),                //                                      .chipselect
		.IO_Pio_avalon_parallel_port_slave_address        (mm_interconnect_0_io_pio_avalon_parallel_port_slave_address),        //     IO_Pio_avalon_parallel_port_slave.address
		.IO_Pio_avalon_parallel_port_slave_write          (mm_interconnect_0_io_pio_avalon_parallel_port_slave_write),          //                                      .write
		.IO_Pio_avalon_parallel_port_slave_read           (mm_interconnect_0_io_pio_avalon_parallel_port_slave_read),           //                                      .read
		.IO_Pio_avalon_parallel_port_slave_readdata       (mm_interconnect_0_io_pio_avalon_parallel_port_slave_readdata),       //                                      .readdata
		.IO_Pio_avalon_parallel_port_slave_writedata      (mm_interconnect_0_io_pio_avalon_parallel_port_slave_writedata),      //                                      .writedata
		.IO_Pio_avalon_parallel_port_slave_byteenable     (mm_interconnect_0_io_pio_avalon_parallel_port_slave_byteenable),     //                                      .byteenable
		.IO_Pio_avalon_parallel_port_slave_chipselect     (mm_interconnect_0_io_pio_avalon_parallel_port_slave_chipselect),     //                                      .chipselect
		.jtag_avalon_jtag_slave_address                   (mm_interconnect_0_jtag_avalon_jtag_slave_address),                   //                jtag_avalon_jtag_slave.address
		.jtag_avalon_jtag_slave_write                     (mm_interconnect_0_jtag_avalon_jtag_slave_write),                     //                                      .write
		.jtag_avalon_jtag_slave_read                      (mm_interconnect_0_jtag_avalon_jtag_slave_read),                      //                                      .read
		.jtag_avalon_jtag_slave_readdata                  (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),                  //                                      .readdata
		.jtag_avalon_jtag_slave_writedata                 (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),                 //                                      .writedata
		.jtag_avalon_jtag_slave_waitrequest               (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest),               //                                      .waitrequest
		.jtag_avalon_jtag_slave_chipselect                (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),                //                                      .chipselect
		.LED_Pio_avalon_parallel_port_slave_address       (mm_interconnect_0_led_pio_avalon_parallel_port_slave_address),       //    LED_Pio_avalon_parallel_port_slave.address
		.LED_Pio_avalon_parallel_port_slave_write         (mm_interconnect_0_led_pio_avalon_parallel_port_slave_write),         //                                      .write
		.LED_Pio_avalon_parallel_port_slave_read          (mm_interconnect_0_led_pio_avalon_parallel_port_slave_read),          //                                      .read
		.LED_Pio_avalon_parallel_port_slave_readdata      (mm_interconnect_0_led_pio_avalon_parallel_port_slave_readdata),      //                                      .readdata
		.LED_Pio_avalon_parallel_port_slave_writedata     (mm_interconnect_0_led_pio_avalon_parallel_port_slave_writedata),     //                                      .writedata
		.LED_Pio_avalon_parallel_port_slave_byteenable    (mm_interconnect_0_led_pio_avalon_parallel_port_slave_byteenable),    //                                      .byteenable
		.LED_Pio_avalon_parallel_port_slave_chipselect    (mm_interconnect_0_led_pio_avalon_parallel_port_slave_chipselect),    //                                      .chipselect
		.sdram_s1_address                                 (mm_interconnect_0_sdram_s1_address),                                 //                              sdram_s1.address
		.sdram_s1_write                                   (mm_interconnect_0_sdram_s1_write),                                   //                                      .write
		.sdram_s1_read                                    (mm_interconnect_0_sdram_s1_read),                                    //                                      .read
		.sdram_s1_readdata                                (mm_interconnect_0_sdram_s1_readdata),                                //                                      .readdata
		.sdram_s1_writedata                               (mm_interconnect_0_sdram_s1_writedata),                               //                                      .writedata
		.sdram_s1_byteenable                              (mm_interconnect_0_sdram_s1_byteenable),                              //                                      .byteenable
		.sdram_s1_readdatavalid                           (mm_interconnect_0_sdram_s1_readdatavalid),                           //                                      .readdatavalid
		.sdram_s1_waitrequest                             (mm_interconnect_0_sdram_s1_waitrequest),                             //                                      .waitrequest
		.sdram_s1_chipselect                              (mm_interconnect_0_sdram_s1_chipselect),                              //                                      .chipselect
		.Switch_Pio_avalon_parallel_port_slave_address    (mm_interconnect_0_switch_pio_avalon_parallel_port_slave_address),    // Switch_Pio_avalon_parallel_port_slave.address
		.Switch_Pio_avalon_parallel_port_slave_write      (mm_interconnect_0_switch_pio_avalon_parallel_port_slave_write),      //                                      .write
		.Switch_Pio_avalon_parallel_port_slave_read       (mm_interconnect_0_switch_pio_avalon_parallel_port_slave_read),       //                                      .read
		.Switch_Pio_avalon_parallel_port_slave_readdata   (mm_interconnect_0_switch_pio_avalon_parallel_port_slave_readdata),   //                                      .readdata
		.Switch_Pio_avalon_parallel_port_slave_writedata  (mm_interconnect_0_switch_pio_avalon_parallel_port_slave_writedata),  //                                      .writedata
		.Switch_Pio_avalon_parallel_port_slave_byteenable (mm_interconnect_0_switch_pio_avalon_parallel_port_slave_byteenable), //                                      .byteenable
		.Switch_Pio_avalon_parallel_port_slave_chipselect (mm_interconnect_0_switch_pio_avalon_parallel_port_slave_chipselect), //                                      .chipselect
		.sys_clk_timer_s1_address                         (mm_interconnect_0_sys_clk_timer_s1_address),                         //                      sys_clk_timer_s1.address
		.sys_clk_timer_s1_write                           (mm_interconnect_0_sys_clk_timer_s1_write),                           //                                      .write
		.sys_clk_timer_s1_readdata                        (mm_interconnect_0_sys_clk_timer_s1_readdata),                        //                                      .readdata
		.sys_clk_timer_s1_writedata                       (mm_interconnect_0_sys_clk_timer_s1_writedata),                       //                                      .writedata
		.sys_clk_timer_s1_chipselect                      (mm_interconnect_0_sys_clk_timer_s1_chipselect),                      //                                      .chipselect
		.sys_id_control_slave_address                     (mm_interconnect_0_sys_id_control_slave_address),                     //                  sys_id_control_slave.address
		.sys_id_control_slave_readdata                    (mm_interconnect_0_sys_id_control_slave_readdata),                    //                                      .readdata
		.sys_pll_pll_slave_address                        (mm_interconnect_0_sys_pll_pll_slave_address),                        //                     sys_pll_pll_slave.address
		.sys_pll_pll_slave_write                          (mm_interconnect_0_sys_pll_pll_slave_write),                          //                                      .write
		.sys_pll_pll_slave_read                           (mm_interconnect_0_sys_pll_pll_slave_read),                           //                                      .read
		.sys_pll_pll_slave_readdata                       (mm_interconnect_0_sys_pll_pll_slave_readdata),                       //                                      .readdata
		.sys_pll_pll_slave_writedata                      (mm_interconnect_0_sys_pll_pll_slave_writedata),                      //                                      .writedata
		.uart_s1_address                                  (mm_interconnect_0_uart_s1_address),                                  //                               uart_s1.address
		.uart_s1_write                                    (mm_interconnect_0_uart_s1_write),                                    //                                      .write
		.uart_s1_read                                     (mm_interconnect_0_uart_s1_read),                                     //                                      .read
		.uart_s1_readdata                                 (mm_interconnect_0_uart_s1_readdata),                                 //                                      .readdata
		.uart_s1_writedata                                (mm_interconnect_0_uart_s1_writedata),                                //                                      .writedata
		.uart_s1_begintransfer                            (mm_interconnect_0_uart_s1_begintransfer),                            //                                      .begintransfer
		.uart_s1_chipselect                               (mm_interconnect_0_uart_s1_chipselect)                                //                                      .chipselect
	);

	niosII_irq_mapper irq_mapper (
		.clk           (sys_pll_c0_clk),                 //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (sys_pll_c0_clk),                     //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (sys_pll_c0_clk),                     //       receiver_clk.clk
		.sender_clk     (sys_pll_c0_clk),                     //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (sys_pll_c0_clk),                     //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),          // reset_in1.reset
		.clk            (sys_pll_c0_clk),                         //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
